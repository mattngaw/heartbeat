`include "./array.sv"

module Testbench;

endmodule: Testbench
